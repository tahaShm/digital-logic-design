library verilog;
use verilog.vl_types.all;
entity testQ4 is
end testQ4;
