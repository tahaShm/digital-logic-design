library verilog;
use verilog.vl_types.all;
entity q7TB is
end q7TB;
