library verilog;
use verilog.vl_types.all;
entity q6TB is
end q6TB;
