library verilog;
use verilog.vl_types.all;
entity testQ2_4 is
end testQ2_4;
