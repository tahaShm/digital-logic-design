library verilog;
use verilog.vl_types.all;
entity counterTB is
end counterTB;
