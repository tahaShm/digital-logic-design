library verilog;
use verilog.vl_types.all;
entity q3TB is
end q3TB;
