library verilog;
use verilog.vl_types.all;
entity testQ2 is
end testQ2;
