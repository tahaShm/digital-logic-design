library verilog;
use verilog.vl_types.all;
entity q14TB is
end q14TB;
