library verilog;
use verilog.vl_types.all;
entity freqTB is
end freqTB;
