library verilog;
use verilog.vl_types.all;
entity q1TB is
end q1TB;
