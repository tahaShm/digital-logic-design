library verilog;
use verilog.vl_types.all;
entity q11TB is
end q11TB;
