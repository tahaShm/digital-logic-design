library verilog;
use verilog.vl_types.all;
entity shiftTB is
end shiftTB;
