library verilog;
use verilog.vl_types.all;
entity testQ1 is
end testQ1;
