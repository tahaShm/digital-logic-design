library verilog;
use verilog.vl_types.all;
entity oc15 is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        d               : in     vl_logic;
        e               : in     vl_logic;
        f               : in     vl_logic;
        g               : in     vl_logic;
        h               : in     vl_logic;
        i               : in     vl_logic;
        j               : in     vl_logic;
        k               : in     vl_logic;
        l               : in     vl_logic;
        m               : in     vl_logic;
        n               : in     vl_logic;
        o               : in     vl_logic;
        y0              : out    vl_logic;
        y1              : out    vl_logic;
        y2              : out    vl_logic;
        y3              : out    vl_logic
    );
end oc15;
