library verilog;
use verilog.vl_types.all;
entity q13TB is
end q13TB;
