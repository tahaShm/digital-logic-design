library verilog;
use verilog.vl_types.all;
entity q4TB is
end q4TB;
