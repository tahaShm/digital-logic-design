library verilog;
use verilog.vl_types.all;
entity q2TB is
end q2TB;
